`timescale 1ns/1ns
module tb_decode5to32();
  reg [4:0] A;
  reg en;
  wire [31:0] out;
  initial begin
    A = 0;
    en = 1;
    #100;
    A = 5'd1;
    #100;
    A = 5'd2;
    #100;
    A = 5'd3;
    #100;
    A = 5'd4;
    #100;
    A = 5'd5;
    #100;
    A = 5'd6;
    #100;
    A = 5'd7;
    #100;
    A = 5'd8;
    #100;
    A = 5'd9;
    #100;
    A = 5'd10;
    #100;
    A = 5'd11;
    #100;
    A = 5'd12;
    #100;
    A = 5'd13;
    #100;
    A = 5'd14;
    #100;
    A = 5'd15;
    #100;
    A = 5'd16;
    #100;
    A = 5'd17;
    #100;
    A = 5'd18;
    #100;
    A = 5'd19;
    #100;
    A = 5'd20;
    #100;
    A = 5'd21;
    #100;
    A = 5'd22;
    #100;
    A = 5'd23;
    #100;
    A = 5'd24;
    #100;
    A = 5'd25;
    #100;
    A = 5'd26;
    #100;
    A = 5'd27;
    #100;
    A = 5'd28;
    #100;
    A = 5'd29;
    #100;
    A = 5'd30;
    #100;
    A = 5'd31;
    #100;
  end
  decode5to32 ins5(
  .A(A),
  .en(en),
  .out(out)
  );
endmodule
    

